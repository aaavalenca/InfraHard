module SignExtend(instruction15_0, instruction31_0);

    input [15:0] instruction15_0;
	output reg[31:0] instruction31_0;

always@(*)
	
	instruction31_0[31:0] = (instruction15_0[15] == 0) ? (32'b00000000000000000000000000000000 + instruction15_0) : (32'b11111111111111110000000000000000 + instruction15_0);

endmodule