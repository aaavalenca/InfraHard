module ShiftLeft2(instructionIn31_0, instructionOut31_0);

    input [31:0] instructionIn31_0;
	output reg [31:0] instructionOut31_0;

always@(*)
	begin
		instructionOut31_0[31:2] = instructionIn31_0[29:0];
		instructionOut31_0[1:0] = 2'b00;
	end
endmodule